module mux_memtoreg(in1, in2 , PC_4 , b , sel , out);
input [31:0] in1, in2 ,PC_4 , b ;
input [1:0] sel;
output reg [31:0]  out ;
//assign #5  PC_4 = 5'b11111 ;
assign #5 b = 5'bxxxxx ;
always @ (in1, in2, PC_4 ,sel)
begin 
case(sel)  
2'b01 : #5 out = in1 ;
2'b00 : #5 out = in2 ;
2'b10 : #5 out = PC_4 ;
2'b11 : #5 out = b ; 
endcase
end 
endmodule 
